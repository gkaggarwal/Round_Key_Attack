-- Written by Gaurav Aggarwal
-- Date: 19th March, 2020
-- Version: v.1.0


LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY Sbox_slice IS
		PORT (SBox_slice_in : IN std_logic_vector (7 downto 0);
		SBox_slice_out : OUT std_logic_vector (7 downto 0));
END SBox_slice;

ARCHITECTURE SBox_slice_logic OF SBox_slice IS
BEGIN
		PROCESS(SBox_slice_in)
		BEGIN
				CASE SBox_slice_in IS 
						 WHEN		X"00"		 =>		SBox_slice_out<=X"63"; 	   
						 WHEN		X"01"		 =>		SBox_slice_out<=X"7c"; 
						 WHEN		X"02"		 =>		SBox_slice_out<=X"77";	  
						 WHEN		X"03"		 =>		SBox_slice_out<=X"7b";	  
						 WHEN		X"04"		 =>		SBox_slice_out<=X"f2";	  
						 WHEN		X"05"		 =>		SBox_slice_out<=X"6b";	  
						 WHEN		X"06"		 =>		SBox_slice_out<=X"6f";	  
						 WHEN		X"07"		 =>		SBox_slice_out<=X"c5";	  
						 WHEN		X"08"		 =>		SBox_slice_out<=X"30";	  
						 WHEN		X"09"		 =>		SBox_slice_out<=X"01";	  
						 WHEN		X"0a"		 =>		SBox_slice_out<=X"67";	  
						 WHEN		X"0b"		 =>		SBox_slice_out<=X"2b";	  
						 WHEN		X"0c"		 =>		SBox_slice_out<=X"fe";	  
						 WHEN		X"0d"		 =>		SBox_slice_out<=X"d7";	  
						 WHEN		X"0e"		 =>		SBox_slice_out<=X"ab";	  
						 WHEN		X"0f"		 =>		SBox_slice_out<=X"76";	  
						 WHEN		X"10"		 =>		SBox_slice_out<=X"ca";	  
						 WHEN		X"11"		 =>		SBox_slice_out<=X"82";	  
						 WHEN		X"12"		 =>		SBox_slice_out<=X"c9";	  
						 WHEN		X"13"		 =>		SBox_slice_out<=X"7d";	  
						 WHEN		X"14"		 =>		SBox_slice_out<=X"fa";	  
						 WHEN		X"15"		 =>		SBox_slice_out<=X"59";	  
						 WHEN		X"16"		 =>		SBox_slice_out<=X"47";	  
						 WHEN		X"17"		 =>		SBox_slice_out<=X"f0";	  
						 WHEN		X"18"		 =>		SBox_slice_out<=X"ad";	  
						 WHEN		X"19"		 =>		SBox_slice_out<=X"d4";	  
						 WHEN		X"1a"		 =>		SBox_slice_out<=X"a2";	  
						 WHEN		X"1b"		 =>		SBox_slice_out<=X"af";	  
						 WHEN		X"1c"		 =>		SBox_slice_out<=X"9c";	  
						 WHEN		X"1d"		 =>		SBox_slice_out<=X"a4";	  
						 WHEN		X"1e"		 =>		SBox_slice_out<=X"72";	  
						 WHEN		X"1f"		 =>		SBox_slice_out<=X"c0";	  
						 WHEN		X"20"		 =>		SBox_slice_out<=X"b7";	  
						 WHEN		X"21"		 =>		SBox_slice_out<=X"fd";	  
						 WHEN		X"22"		 =>		SBox_slice_out<=X"93";	  
						 WHEN		X"23"		 =>		SBox_slice_out<=X"26";	  
						 WHEN		X"24"		 =>		SBox_slice_out<=X"36";	  
						 WHEN		X"25"		 =>		SBox_slice_out<=X"3f";	  
						 WHEN		X"26"		 =>		SBox_slice_out<=X"f7";	  
						 WHEN		X"27"		 =>		SBox_slice_out<=X"cc";	  
						 WHEN		X"28"		 =>		SBox_slice_out<=X"34";	  
						 WHEN		X"29"		 =>		SBox_slice_out<=X"a5";	  
						 WHEN		X"2a"		 =>		SBox_slice_out<=X"e5";	  
						 WHEN		X"2b"		 =>		SBox_slice_out<=X"f1";	  
						 WHEN		X"2c"		 =>		SBox_slice_out<=X"71";	  
						 WHEN		X"2d"		 =>		SBox_slice_out<=X"d8";	  
						 WHEN		X"2e"		 =>		SBox_slice_out<=X"31";	  
						 WHEN		X"2f"		 =>		SBox_slice_out<=X"15";	  
						 WHEN		X"30"		 =>		SBox_slice_out<=X"04";	  
						 WHEN		X"31"		 =>		SBox_slice_out<=X"c7";	  
						 WHEN		X"32"		 =>		SBox_slice_out<=X"23";	  
						 WHEN		X"33"		 =>		SBox_slice_out<=X"c3";	  
						 WHEN		X"34"		 =>		SBox_slice_out<=X"18";	  
						 WHEN		X"35"		 =>		SBox_slice_out<=X"96";	  
						 WHEN		X"36"		 =>		SBox_slice_out<=X"05";	  
						 WHEN		X"37"		 =>		SBox_slice_out<=X"9a";	  
						 WHEN		X"38"		 =>		SBox_slice_out<=X"07";	  
						 WHEN		X"39"		 =>		SBox_slice_out<=X"12";	  
						 WHEN		X"3a"		 =>		SBox_slice_out<=X"80";	  
						 WHEN		X"3b"		 =>		SBox_slice_out<=X"e2";	  
						 WHEN		X"3c"		 =>		SBox_slice_out<=X"eb";	  
						 WHEN		X"3d"		 =>		SBox_slice_out<=X"27";	  
						 WHEN		X"3e"		 =>		SBox_slice_out<=X"b2";	  
						 WHEN		X"3f"		 =>		SBox_slice_out<=X"75";	  
						 WHEN		X"40"		 =>		SBox_slice_out<=X"09";	  
						 WHEN		X"41"		 =>		SBox_slice_out<=X"83";	  
						 WHEN		X"42"		 =>		SBox_slice_out<=X"2c";	  
						 WHEN		X"43"		 =>		SBox_slice_out<=X"1a";	  
						 WHEN		X"44"		 =>		SBox_slice_out<=X"1b";	  
						 WHEN		X"45"		 =>		SBox_slice_out<=X"6e";	  
						 WHEN		X"46"		 =>		SBox_slice_out<=X"5a";	  
						 WHEN		X"47"		 =>		SBox_slice_out<=X"a0";	  
						 WHEN		X"48"		 =>		SBox_slice_out<=X"52";	  
						 WHEN		X"49"		 =>		SBox_slice_out<=X"3b";	  
						 WHEN		X"4a"		 =>		SBox_slice_out<=X"d6";	  
						 WHEN		X"4b"		 =>		SBox_slice_out<=X"b3";	  
						 WHEN		X"4c"		 =>		SBox_slice_out<=X"29";	  
						 WHEN		X"4d"		 =>		SBox_slice_out<=X"e3";	  
						 WHEN		X"4e"		 =>		SBox_slice_out<=X"2f";	  
						 WHEN		X"4f"		 =>		SBox_slice_out<=X"84";	  
						 WHEN		X"50"		 =>		SBox_slice_out<=X"53";	  
						 WHEN		X"51"		 =>		SBox_slice_out<=X"d1";	  
						 WHEN		X"52"		 =>		SBox_slice_out<=X"00";	  
						 WHEN		X"53"		 =>		SBox_slice_out<=X"ed";	  
						 WHEN		X"54"		 =>		SBox_slice_out<=X"20";	  
						 WHEN		X"55"		 =>		SBox_slice_out<=X"fc";	  
						 WHEN		X"56"		 =>		SBox_slice_out<=X"b1";	  
						 WHEN		X"57"		 =>		SBox_slice_out<=X"5b";	  
						 WHEN		X"58"		 =>		SBox_slice_out<=X"6a";	  
						 WHEN		X"59"		 =>		SBox_slice_out<=X"cb";	  
						 WHEN		X"5a"		 =>		SBox_slice_out<=X"be";	  
						 WHEN		X"5b"		 =>		SBox_slice_out<=X"39";	  
						 WHEN		X"5c"		 =>		SBox_slice_out<=X"4a";	  
						 WHEN		X"5d"		 =>		SBox_slice_out<=X"4c";	  
						 WHEN		X"5e"		 =>		SBox_slice_out<=X"58";	  
						 WHEN		X"5f"		 =>		SBox_slice_out<=X"cf";	  
						 WHEN		X"60"		 =>		SBox_slice_out<=X"d0";	  
						 WHEN		X"61"		 =>		SBox_slice_out<=X"ef";	  
						 WHEN		X"62"		 =>		SBox_slice_out<=X"aa";	  
						 WHEN		X"63"		 =>		SBox_slice_out<=X"fb";	  
						 WHEN		X"64"		 =>		SBox_slice_out<=X"43";	  
						 WHEN		X"65"		 =>		SBox_slice_out<=X"4d";	  
						 WHEN		X"66"		 =>		SBox_slice_out<=X"33";	  
						 WHEN		X"67"		 =>		SBox_slice_out<=X"85";	  
						 WHEN		X"68"		 =>		SBox_slice_out<=X"45";	  
						 WHEN		X"69"		 =>		SBox_slice_out<=X"f9";	  
						 WHEN		X"6a"		 =>		SBox_slice_out<=X"02";	  
						 WHEN		X"6b"		 =>		SBox_slice_out<=X"7f";	  
						 WHEN		X"6c"		 =>		SBox_slice_out<=X"50";	  
						 WHEN		X"6d"		 =>		SBox_slice_out<=X"3c";	  
						 WHEN		X"6e"		 =>		SBox_slice_out<=X"9f";	  
						 WHEN		X"6f"		 =>		SBox_slice_out<=X"a8";	  
						 WHEN		X"70"		 =>		SBox_slice_out<=X"51";	  
						 WHEN		X"71"		 =>		SBox_slice_out<=X"a3";	  
						 WHEN		X"72"		 =>		SBox_slice_out<=X"40";	  
						 WHEN		X"73"		 =>		SBox_slice_out<=X"8f";	  
						 WHEN		X"74"		 =>		SBox_slice_out<=X"92";	  
						 WHEN		X"75"		 =>		SBox_slice_out<=X"9d";	  
						 WHEN		X"76"		 =>		SBox_slice_out<=X"38";	  
						 WHEN		X"77"		 =>		SBox_slice_out<=X"f5";	  
						 WHEN		X"78"		 =>		SBox_slice_out<=X"bc";	  
						 WHEN		X"79"		 =>		SBox_slice_out<=X"b6";	  
						 WHEN		X"7a"		 =>		SBox_slice_out<=X"da";	  
						 WHEN		X"7b"		 =>		SBox_slice_out<=X"21";	  
						 WHEN		X"7c"		 =>		SBox_slice_out<=X"10";	  
						 WHEN		X"7d"		 =>		SBox_slice_out<=X"ff";	  
						 WHEN		X"7e"		 =>		SBox_slice_out<=X"f3";	  
						 WHEN		X"7f"		 =>		SBox_slice_out<=X"d2";	  
						 WHEN		X"80"		 =>		SBox_slice_out<=X"cd";	  
						 WHEN		X"81"		 =>		SBox_slice_out<=X"0c";	  
						 WHEN		X"82"		 =>		SBox_slice_out<=X"13";	  
						 WHEN		X"83"		 =>		SBox_slice_out<=X"ec";	  
						 WHEN		X"84"		 =>		SBox_slice_out<=X"5f";	  
						 WHEN		X"85"		 =>		SBox_slice_out<=X"97";	  
						 WHEN		X"86"		 =>		SBox_slice_out<=X"44";	  
						 WHEN		X"87"		 =>		SBox_slice_out<=X"17";	  
						 WHEN		X"88"		 =>		SBox_slice_out<=X"c4";	  
						 WHEN		X"89"		 =>		SBox_slice_out<=X"a7";	  
						 WHEN		X"8a"		 =>		SBox_slice_out<=X"7e";	  
						 WHEN		X"8b"		 =>		SBox_slice_out<=X"3d";	  
						 WHEN		X"8c"		 =>		SBox_slice_out<=X"64";	  
						 WHEN		X"8d"		 =>		SBox_slice_out<=X"5d";	  
						 WHEN		X"8e"		 =>		SBox_slice_out<=X"19";	  
						 WHEN		X"8f"		 =>		SBox_slice_out<=X"73";	  
						 WHEN		X"90"		 =>		SBox_slice_out<=X"60";	  
						 WHEN		X"91"		 =>		SBox_slice_out<=X"81";	  
						 WHEN		X"92"		 =>		SBox_slice_out<=X"4f";	  
						 WHEN		X"93"		 =>		SBox_slice_out<=X"dc";	  
						 WHEN		X"94"		 =>		SBox_slice_out<=X"22";	  
						 WHEN		X"95"		 =>		SBox_slice_out<=X"2a";	  
						 WHEN		X"96"		 =>		SBox_slice_out<=X"90";	  
						 WHEN		X"97"		 =>		SBox_slice_out<=X"88";	  
						 WHEN		X"98"		 =>		SBox_slice_out<=X"46";	  
						 WHEN		X"99"		 =>		SBox_slice_out<=X"ee";	  
						 WHEN		X"9a"		 =>		SBox_slice_out<=X"b8";	  
						 WHEN		X"9b"		 =>		SBox_slice_out<=X"14";	  
						 WHEN		X"9c"		 =>		SBox_slice_out<=X"de";	  
						 WHEN		X"9d"		 =>		SBox_slice_out<=X"5e";	  
						 WHEN		X"9e"		 =>		SBox_slice_out<=X"0b";	  
						 WHEN		X"9f"		 =>		SBox_slice_out<=X"db";	  
						 WHEN		X"a0"		 =>		SBox_slice_out<=X"e0";	  
						 WHEN		X"a1"		 =>		SBox_slice_out<=X"32";	  
						 WHEN		X"a2"		 =>		SBox_slice_out<=X"3a";	  
						 WHEN		X"a3"		 =>		SBox_slice_out<=X"0a";	  
						 WHEN		X"a4"		 =>		SBox_slice_out<=X"49";	  
						 WHEN		X"a5"		 =>		SBox_slice_out<=X"06";	  
						 WHEN		X"a6"		 =>		SBox_slice_out<=X"24";	  
						 WHEN		X"a7"		 =>		SBox_slice_out<=X"5c";	  
						 WHEN		X"a8"		 =>		SBox_slice_out<=X"c2";	  
						 WHEN		X"a9"		 =>		SBox_slice_out<=X"d3";	  
						 WHEN		X"aa"		 =>		SBox_slice_out<=X"ac";	  
						 WHEN		X"ab"		 =>		SBox_slice_out<=X"62";	  
						 WHEN		X"ac"		 =>		SBox_slice_out<=X"91";	  
						 WHEN		X"ad"		 =>		SBox_slice_out<=X"95";	  
						 WHEN		X"ae"		 =>		SBox_slice_out<=X"e4";	  
						 WHEN		X"af"		 =>		SBox_slice_out<=X"79";	  
						 WHEN		X"b0"		 =>		SBox_slice_out<=X"e7";	  
						 WHEN		X"b1"		 =>		SBox_slice_out<=X"c8";	  
						 WHEN		X"b2"		 =>		SBox_slice_out<=X"37";	  
						 WHEN		X"b3"		 =>		SBox_slice_out<=X"6d";	  
						 WHEN		X"b4"		 =>		SBox_slice_out<=X"8d";	  
						 WHEN		X"b5"		 =>		SBox_slice_out<=X"d5";	  
						 WHEN		X"b6"		 =>		SBox_slice_out<=X"4e";	  
						 WHEN		X"b7"		 =>		SBox_slice_out<=X"a9";	  
						 WHEN		X"b8"		 =>		SBox_slice_out<=X"6c";	  
						 WHEN		X"b9"		 =>		SBox_slice_out<=X"56";	  
						 WHEN		X"ba"		 =>		SBox_slice_out<=X"f4";	  
						 WHEN		X"bb"		 =>		SBox_slice_out<=X"ea";	  
						 WHEN		X"bc"		 =>		SBox_slice_out<=X"65";	  
						 WHEN		X"bd"		 =>		SBox_slice_out<=X"7a";	  
						 WHEN		X"be"		 =>		SBox_slice_out<=X"ae";	  
						 WHEN		X"bf"		 =>		SBox_slice_out<=X"08";	  
						 WHEN		X"c0"		 =>		SBox_slice_out<=X"ba";	  
						 WHEN		X"c1"		 =>		SBox_slice_out<=X"78";	  
						 WHEN		X"c2"		 =>		SBox_slice_out<=X"25";	  
						 WHEN		X"c3"		 =>		SBox_slice_out<=X"2e";	  
						 WHEN		X"c4"		 =>		SBox_slice_out<=X"1c";	  
						 WHEN		X"c5"		 =>		SBox_slice_out<=X"a6";	  
						 WHEN		X"c6"		 =>		SBox_slice_out<=X"b4";	  
						 WHEN		X"c7"		 =>		SBox_slice_out<=X"c6";	  
						 WHEN		X"c8"		 =>		SBox_slice_out<=X"e8";	  
						 WHEN		X"c9"		 =>		SBox_slice_out<=X"dd";	  
						 WHEN		X"ca"		 =>		SBox_slice_out<=X"74";	  
						 WHEN		X"cb"		 =>		SBox_slice_out<=X"1f";	  
						 WHEN		X"cc"		 =>		SBox_slice_out<=X"4b";	  
						 WHEN		X"cd"		 =>		SBox_slice_out<=X"bd";	  
						 WHEN		X"ce"		 =>		SBox_slice_out<=X"8b";	  
						 WHEN		X"cf"		 =>		SBox_slice_out<=X"8a";	  
						 WHEN		X"d0"		 =>		SBox_slice_out<=X"70";	  
						 WHEN		X"d1"		 =>		SBox_slice_out<=X"3e";	  
						 WHEN		X"d2"		 =>		SBox_slice_out<=X"b5";	  
						 WHEN		X"d3"		 =>		SBox_slice_out<=X"66";	  
						 WHEN		X"d4"		 =>		SBox_slice_out<=X"48";	  
						 WHEN		X"d5"		 =>		SBox_slice_out<=X"03";	  
						 WHEN		X"d6"		 =>		SBox_slice_out<=X"f6";	  
						 WHEN		X"d7"		 =>		SBox_slice_out<=X"0e";	  
						 WHEN		X"d8"		 =>		SBox_slice_out<=X"61";	  
						 WHEN		X"d9"		 =>		SBox_slice_out<=X"35";	  
						 WHEN		X"da"		 =>		SBox_slice_out<=X"57";	  
						 WHEN		X"db"		 =>		SBox_slice_out<=X"b9";	  
						 WHEN		X"dc"		 =>		SBox_slice_out<=X"86";	  
						 WHEN		X"dd"		 =>		SBox_slice_out<=X"c1";	  
						 WHEN		X"de"		 =>		SBox_slice_out<=X"1d";	  
						 WHEN		X"df"		 =>		SBox_slice_out<=X"9e";	  
						 WHEN		X"e0"		 =>		SBox_slice_out<=X"e1";	  
						 WHEN		X"e1"		 =>		SBox_slice_out<=X"f8";	  
						 WHEN		X"e2"		 =>		SBox_slice_out<=X"98";	  
						 WHEN		X"e3"		 =>		SBox_slice_out<=X"11";	  
						 WHEN		X"e4"		 =>		SBox_slice_out<=X"69";	  
						 WHEN		X"e5"		 =>		SBox_slice_out<=X"d9";	  
						 WHEN		X"e6"		 =>		SBox_slice_out<=X"8e";	  
						 WHEN		X"e7"		 =>		SBox_slice_out<=X"94";	  
						 WHEN		X"e8"		 =>		SBox_slice_out<=X"9b";	  
						 WHEN		X"e9"		 =>		SBox_slice_out<=X"1e";	  
						 WHEN		X"ea"		 =>		SBox_slice_out<=X"87";	  
						 WHEN		X"eb"		 =>		SBox_slice_out<=X"e9";	  
						 WHEN		X"ec"		 =>		SBox_slice_out<=X"ce";	  
						 WHEN		X"ed"		 =>		SBox_slice_out<=X"55";	  
						 WHEN		X"ee"		 =>		SBox_slice_out<=X"28";	  
						 WHEN		X"ef"		 =>		SBox_slice_out<=X"df";	  
						 WHEN		X"f0"		 =>		SBox_slice_out<=X"8c";	  
						 WHEN		X"f1"		 =>		SBox_slice_out<=X"a1";	  
						 WHEN		X"f2"		 =>		SBox_slice_out<=X"89";	  
						 WHEN		X"f3"		 =>		SBox_slice_out<=X"0d";	  
						 WHEN		X"f4"		 =>		SBox_slice_out<=X"bf";	  
						 WHEN		X"f5"		 =>		SBox_slice_out<=X"e6";	  
						 WHEN		X"f6"		 =>		SBox_slice_out<=X"42";	  
						 WHEN		X"f7"		 =>		SBox_slice_out<=X"68";	  
						 WHEN		X"f8"		 =>		SBox_slice_out<=X"41";	  
						 WHEN		X"f9"		 =>		SBox_slice_out<=X"99";	  
						 WHEN		X"fa"		 =>		SBox_slice_out<=X"2d";	  
						 WHEN		X"fb"		 =>		SBox_slice_out<=X"0f";	  
						 WHEN		X"fc"		 =>		SBox_slice_out<=X"b0";	  
						 WHEN		X"fd"		 =>		SBox_slice_out<=X"54";	  
						 WHEN		X"fe"		 =>		SBox_slice_out<=X"bb";	  
						 WHEN       X"ff"		 =>     SBox_slice_out<=X"16";
						 WHEN others             =>     SBox_slice_out<=X"16";
				 END CASE;
		 END PROCESS;
END SBox_slice_logic;
